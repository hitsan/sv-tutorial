// パイプライン化された乗算器の各種実装 - テストベンチ
// テストベンチは実装ごとに分割しました。
// - multiplier_pipelined_multistage_tb.sv
// - multiplier_pipelined_array_tb.sv

`timescale 1ns / 100ps
