// 演習1: 基本的なモジュールインスタンス化
// 4:1マルチプレクサを2:1マルチプレクサから構成

/*
 * 要求仕様:
 * - 2:1マルチプレクサ3個を使って4:1マルチプレクサを実装
 * - ../combinational/examples/mux2x1.sv を使用
 *
 * 構造:
 *           ┌───────┐
 *    in[0]──┤       │
 *           │ MUX0  ├──┐
 *    in[1]──┤       │  │  ┌───────┐
 *           └───────┘  ├──┤       │
 *    sel[0]────────────┘  │       │
 *                         │ MUX2  ├── out
 *           ┌───────┐  ┌──┤       │
 *    in[2]──┤       │  │  └───────┘
 *           │ MUX1  ├──┘
 *    in[3]──┤       │
 *           └───────┘
 *    sel[0]────────────┘
 *    sel[1]──────────────────────┘
 */

module mux4x1_structural (
    input  logic [3:0] in,
    input  logic [1:0] sel,
    output logic       out
);
    // ここに実装
    // ヒント: mux2x1を3個インスタンス化する

endmodule : mux4x1_structural
