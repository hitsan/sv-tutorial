`timescale 1ns/1ps
module direct_mapped_cache_tb;
    initial begin
        $display("direct_mapped_cache_tb: TODO");
        $finish;
    end
endmodule
