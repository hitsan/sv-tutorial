`timescale 1ns/1ps
module hw_scheduler_tb;
    initial begin
        $display("hw_scheduler_tb: TODO");
        $finish;
    end
endmodule
