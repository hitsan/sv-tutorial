`timescale 1ns/1ps
module dma_m2s_tb;
    initial begin
        $display("dma_m2s_tb: TODO");
        $finish;
    end
endmodule
