`timescale 1ns/1ps
module eth_rx_parser_tb;
    // TODO: テストベンチ実装
    initial begin
        $display("eth_rx_parser_tb: TODO - Implementation pending");
        $finish;
    end
endmodule
