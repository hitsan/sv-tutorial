// パイプライン化された乗算器の各種実装
// 2つの実装を別ファイルに分割しました。
// - multiplier_pipelined_multistage.sv
// - multiplier_pipelined_array.sv

`timescale 1ns / 100ps
