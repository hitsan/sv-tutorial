// priority_encoder_4in のテストベンチ
// 全16パターンを網羅的にテストし、assertionでエラーを検出

`timescale 1ns / 100ps

module priority_encoder_4in_tb;

    // ============================================================================
    // テストベンチの信号宣言
    // ============================================================================
    logic [3:0] data_in;
    logic [1:0] data_out;

    // ============================================================================
    // DUT (Device Under Test) のインスタンス化
    // ============================================================================
    priority_encoder_4in DUT (.*);

    // ============================================================================
    // Golden Reference関数
    // ============================================================================
    // DUTの期待値を計算する関数
    // 最上位ビットから優先的にエンコード
    function automatic logic [1:0] calc_expected(logic [3:0] din);
        if (din[3]) return 2'b11;
        else if (din[2]) return 2'b10;
        else if (din[1]) return 2'b01;
        else return 2'b00;  // din[0]=1 or all 0
    endfunction

    // ============================================================================
    // テストケース実行タスク
    // ============================================================================
    task automatic test_case(input logic [3:0] din);
        logic [1:0] expected;

        // 入力を設定
        data_in = din;

        // 組み合わせ回路なので伝搬遅延を考慮
        #1;

        // 期待値を計算
        expected = calc_expected(din);

        // 出力が期待値と一致することを確認（===でX/Z値も厳密にチェック）
        assert (data_out === expected)
            else $error("[%0t] data_in=4'b%b: data_out=%b expected=%b",
                        $realtime, din, data_out, expected);

        #1;  // 次のテストケースまで待機
    endtask

    // ============================================================================
    // テストシーケンス
    // ============================================================================
    initial begin
        // 時刻フォーマット設定
        $timeformat(-9, 0, " ns");

        // テスト開始メッセージ
        $display("=================================================");
        $display("Priority Encoder 4-input Test");
        $display("=================================================");

        // 全16パターンをテスト（4'b0000 ～ 4'b1111）
        for (int i = 0; i < 16; i++) begin
            test_case(i[3:0]);
        end

        // テスト終了
        $display("=================================================");
        $display("Tests completed.");
        $display("=================================================");
        $finish;
    end

    // ============================================================================
    // タイムアウト保護
    // ============================================================================
    initial begin
        #1000;  // 最大シミュレーション時間
        $display("ERROR: Simulation timeout!");
        $finish;
    end

endmodule : priority_encoder_4in_tb


// ============================================================================
// テストベンチ設計のポイント
// ============================================================================
// 1. 全16パターンを網羅的にテスト（完全なカバレッジ）
// 2. Golden reference関数で期待値を自動計算
// 3. assertを使って自動的にエラーを検出
// 4. === 演算子でX/Z値も厳密にチェック
// 5. タイムアウト保護でハングを防ぐ
// 6. ブロッキング代入 (=) を使用（組み合わせ回路）
//
// 動作確認:
// - エラーなしで "Tests completed." が表示されることを確認
// - エラー時は該当の入力値と期待値/実際値が表示される
