// パイプライン化された乗算器の各種実装
// 様々なアーキテクチャのパイプライン乗算器を学習するための実装集
//
// このファイルには5つの異なるパイプラインアーキテクチャが含まれています:
// 1. Multi-Stage Pipeline: 基本的な3ステージパイプライン
// 2. Booth Encoding: Radix-2 Booth符号化による部分積削減
// 3. Wallace Tree: 並列加算ツリーによる高速化
// 4. Array Multiplier: シストリックアレイ構造
// 5. Carry-Save: キャリーセーブ演算による規則的削減

`timescale 1ns / 100ps

// ============================================================================
// 例1: Multi-Stage Pipeline (3ステージ)
// ============================================================================
// 要件:
// - 基本的な2ステージパイプラインを3ステージに拡張
// - 各ステージでバランスよく処理を分散
//
// 学習ポイント:
// - パイプラインステージ数とレイテンシの関係
// - ステージ数を増やすことでクリティカルパスを短縮
// - レイテンシは増加するがスループットは維持
//
// パイプライン構成:
// - Stage 1: 入力レジスタ (in0_r, in1_r)
// - Stage 2: 乗算レジスタ (mul_r)
// - Stage 3: 出力レジスタ (product)
//
module multiplier_pipelined_multistage #(
    parameter int INPUT_WIDTH = 8,
    localparam int OUTPUT_WIDTH = INPUT_WIDTH * 2
) (
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic [INPUT_WIDTH-1:0]   in0,
    input  logic [INPUT_WIDTH-1:0]   in1,
    output logic [OUTPUT_WIDTH-1:0]  product
);
  logic [INPUT_WIDTH-1:0] in0_r;
  logic [INPUT_WIDTH-1:0] in1_r;
  logic [OUTPUT_WIDTH-1:0] mul_r;
  always_ff @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      in0_r <= '0;
      in1_r <= '0;
      product <= '0;
    end else begin
      in0_r <= in0;
      in1_r <= in1;
      mul_r <= in0_r * in1_r;
      product <= mul_r;
    end
  end
endmodule : multiplier_pipelined_multistage


// ============================================================================
// 例2: Booth Encoding Pipeline (Radix-2)
// ============================================================================
// 要件:
// - Radix-2 Boothアルゴリズムによる部分積削減
// - 3ステージパイプライン: エンコード → 部分積生成 → 累算
// - 符号付き演算を自然に処理
//
// Booth Encoding (Radix-2)の真理値表:
// 乗数のビットペア [i+1, i, i-1] を見て動作を決定
//   000 → 0
//   001 → +multiplicand
//   010 → +multiplicand
//   011 → +2*multiplicand
//   100 → -2*multiplicand
//   101 → -multiplicand
//   110 → -multiplicand
//   111 → 0
//
// 学習ポイント:
// - アルゴリズムによる部分積数の削減（8個→4-5個）
// - 符号付き演算がハードウェアで自然に処理される仕組み
// - ハードウェアとアルゴリズムの関係
// - Boothアルゴリズムが特にsigned乗算で有利な理由
//
// 実装ヒント（教育的簡略版）:
// - 完全なBoothアルゴリズムは複雑なため、基本構造のみ実装
// - Stage 1: 入力レジスタ
// - Stage 2: 乗数を1ビット拡張（Booth用）
// - Stage 3: 乗算実行 + 出力
// - IS_SIGNEDでsigned/unsignedを切り替え（generateまたはif文）
//
module multiplier_pipelined_booth #(
    parameter int INPUT_WIDTH = 8,
    parameter bit IS_SIGNED = 1'b1,  // Boothはsignedに有利
    localparam int OUTPUT_WIDTH = INPUT_WIDTH * 2
) (
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic [INPUT_WIDTH-1:0]   in0,
    input  logic [INPUT_WIDTH-1:0]   in1,
    output logic [OUTPUT_WIDTH-1:0]  product
);

    // TODO: Boothエンコーディングを使用した3ステージパイプラインを実装
    // - IS_SIGNEDパラメータでsigned/unsigned乗算を切り替え
    // - signed版ではsigned'()キャストを使用

endmodule : multiplier_pipelined_booth


// ============================================================================
// 例3: Wallace Tree Pipeline
// ============================================================================
// 要件:
// - 部分積を並列に削減するWallace Tree構造
// - 3:2 Compressor (CSA) を使用した削減
// - 4ステージパイプライン: 部分積生成 → 削減層1 → 削減層2 → CPA
//
// Wallace Tree アルゴリズム (8x8):
// - 8個の部分積を生成
// - 3:2 CSAで並列に削減: 8 → 6 → 4 → 2
// - 最終的に2つのベクタ（sum + carry）をCPAで加算
//
// 学習ポイント:
// - 並列削減による高速化
// - 3:2圧縮器（Full Adder）の活用
// - 不規則だが最適化された構造
//
// 実装ヒント:
// - CSA (3:2 Compressor) 関数を定義
//   sum = a ^ b ^ c
//   carry = ((a & b) | (b & c) | (a & c)) << 1
// - Stage 1: 部分積生成 pp[i] = in1[i] ? (in0 << i) : 0
// - Stage 2-3: CSAで段階的に削減
// - Stage 4: 最終加算
//
module multiplier_pipelined_wallace #(
    parameter int INPUT_WIDTH = 8,
    localparam int OUTPUT_WIDTH = INPUT_WIDTH * 2
) (
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic [INPUT_WIDTH-1:0]   in0,
    input  logic [INPUT_WIDTH-1:0]   in1,
    output logic [OUTPUT_WIDTH-1:0]  product
);

    // TODO: Wallace Treeを使用した4ステージパイプラインを実装
    // - 3:2 CSA関数を定義
    // - 部分積を生成
    // - CSAで段階的に削減
    // - 最終的にCPAで加算

endmodule : multiplier_pipelined_wallace


// ============================================================================
// 例4: Array Multiplier Pipeline
// ============================================================================
// 要件:
// - シストリックアレイ構造の乗算器
// - 各行が1パイプラインステージ
// - 規則的で理解しやすい構造
//
// アレイ乗算器:
// - 8x8の2次元配列構造（概念的）
// - 各行: 部分積を生成し、前の行の結果に加算
// - 行ごとにパイプラインレジスタを配置
//
// 学習ポイント:
// - シストリックアレイアーキテクチャ
// - 規則的な構造の利点（設計・検証が容易）
// - 空間パイプライン vs 時間パイプライン
// - レイテンシは長いが、構造が単純
//
// 実装ヒント:
// - 各行でsum/carryレジスタを保持
// - 第i行: 部分積 pp[i] を前の行の結果に加算
// - INPUT_WIDTH個のステージ（8ステージ）
//
module multiplier_pipelined_array #(
    parameter int INPUT_WIDTH = 8,
    localparam int OUTPUT_WIDTH = INPUT_WIDTH * 2
) (
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic [INPUT_WIDTH-1:0]   in0,
    input  logic [INPUT_WIDTH-1:0]   in1,
    output logic [OUTPUT_WIDTH-1:0]  product
);

    // TODO: アレイ乗算器のパイプライン構造を実装
    // - 各行のレジスタを定義（row_sum, row_carry）
    // - 各行で部分積を生成し、前の行の結果に加算
    // - 最終行の結果を出力

endmodule : multiplier_pipelined_array


// ============================================================================
// 例5: Carry-Save Pipeline
// ============================================================================
// 要件:
// - キャリーセーブ演算を使用した規則的削減
// - 中間結果をsum/carry形式で保持
// - 最終段のみキャリー伝搬加算
//
// Carry-Save Algorithm:
// - 3:2 CSAで系統的に削減
// - Wallace Treeより規則的
// - 4ステージ: 部分積生成 → CSA削減1 → CSA削減2 → CPA
//
// 学習ポイント:
// - キャリーセーブ演算の原理
// - 冗長表現（sum + carry）の利点
// - 規則的削減 vs 最適削減のトレードオフ
//
// 実装ヒント:
// - CSA関数を定義（Wallace Treeと同じ）
// - Stage 1: 部分積生成
// - Stage 2-3: CSAで削減（sum/carry分離を維持）
// - Stage 4: 最終CPA
//
module multiplier_pipelined_csa #(
    parameter int INPUT_WIDTH = 8,
    localparam int OUTPUT_WIDTH = INPUT_WIDTH * 2
) (
    input  logic                     clk,
    input  logic                     rst_n,
    input  logic [INPUT_WIDTH-1:0]   in0,
    input  logic [INPUT_WIDTH-1:0]   in1,
    output logic [OUTPUT_WIDTH-1:0]  product
);

    // TODO: Carry-Saveパイプラインを実装
    // - CSA (3:2 Compressor) 関数を定義
    // - 4ステージのパイプライン構造
    // - sum/carry形式を最終段まで保持

endmodule : multiplier_pipelined_csa
