`timescale 1ns/1ps
module udp_tx_tb;
    initial begin
        $display("udp_tx_tb: TODO");
        $finish;
    end
endmodule
