// Greg Stitt
// University of Florida

`timescale 1ns / 100ps

module multiplier_tb;

endmodule
