`timescale 1ns/1ps
module udp_rx_tb;
    initial begin
        $display("udp_rx_tb: TODO");
        $finish;
    end
endmodule
