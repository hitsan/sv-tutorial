`timescale 1ns/1ps
module simple_udp_loopback_tb;
    initial begin
        $display("simple_udp_loopback_tb: TODO");
        $finish;
    end
endmodule
